* TOPOLOGIA 8T-SER

.TITLE '8T-SER 0.5GHz'

.OPTION POST = 2
* .PRINT v(q) v(qb) v(q2) v(q2b) v(bit) v(we) v(wl) v(pre) v(sae)

.include 7nm_TT.pm

.include Leitura.cir
.include Escrita.cir
.include PreCarga.cir

* PARAMETROS
.param fin_auxiliares = 1
.param fin = 1

* TENSAO DO CIRCUITO
.param supply = 0.7

* TEMPOS
.param clock = 0.5g
.param slope = '0.01*period'
.param period = '1/clock'
.param step = 'period/7'

.global supply gnd

* SUPPLY DO CIRCUITO
Vvdd vdd gnd DC supply

* SIMULACAO

Vbit bit gnd PWL(0ns 0 '2*period' 0 '2*period+slope' supply)

Vwe we gnd PWL(0ns supply 'period' supply 'period + slope' 0
+ '2*period' 0 '2*period + slope' supply
+ '3*period' supply '3*period + slope' 0)

Vwl wl gnd PWL(0ns 0 '3*step' 0 '3*step + slope' supply '4*step' supply '4*step + slope' 0
+ 'period + 3*step' 0 'period + 3*step + slope' supply 'period + 4*step' supply 'period + 4*step + slope' 0
+ '2*period + 3*step' 0 '2*period + 3*step + slope' supply '2*period + 4*step' supply '2*period + 4*step + slope' 0
+ '3*period + 3*step' 0 '3*period + 3*step + slope' supply '3*period + 4*step' supply '3*period + 4*step + slope' 0)

Vpre 	pre	    gnd		PWL ( '0*step'              supply  'step'                supply
+ 'step+slope'          0       '6*step'              0
+ '6*step+slope'        supply  'period+step'           supply
+ 'period+step+slope'     0       'period+6*step'         0
+ 'period+6*step+slope'   supply  '2*period+step'		  supply
+ '2*period+step+slope'   0       '2*period+6*step'       0
+ '2*period+6*step+slope' supply  '3*period+step'         supply
+ '3*period+step+slope'   0       '3*period+6*step'       0
+ '3*period+6*step+slope' supply  '4*period'		      supply)

Vsae 	sae	    gnd		PWL ( '0*step'              supply  'period+4*step'         supply
+ 'period+4*step+slope'   0       'period+5*step'         0
+ 'period+5*step+slope'   supply  '3*period+4*step'       supply
+ '3*period+4*step+slope' 0       '3*period+5*step'       0
+ '3*period+5*step+slope' supply  '4*period'              supply)


* DECLARACAO DO CIRCUITO

*  CIRCUITOS AUXILIARES

* PRE-CARGA
Xprecarga pre bl blb vdd gnd pre_carga fin=fin_auxiliares

* ESCRITA
Xescrita  bit we bl blb vdd gnd escrita fin=fin_auxiliares

* LEITURA
Xleitura sae bl blb out outb vdd gnd leitura fin=fin_auxiliares

* CELULA

*Pull-UP
Mp1     vdd     q2      qb     vdd   pmos_rvt   nfin = fin
Mp2     q         q2b     vdd  vdd   pmos_rvt   nfin = fin
Mp3     vdd     q2b     q2     vdd   pmos_rvt   nfin = fin
Mp4     q2b       q2      vdd  vdd   pmos_rvt   nfin = fin

*Access WL
Mn1     wl        q       qb     gnd     nmos_rvt   nfin = fin
Mn2     q         qb      wl     gnd     nmos_rvt   nfin = fin

*Access Bitlines
Mn3     bl        qb      q2     gnd     nmos_rvt   nfin = fin
Mn4     q2b       q       blb    gnd     nmos_rvt   nfin = fin


* CAPACITORES
Cload	out gnd	1f
Cload2	outb gnd 1f


* VALOR INICIAL DA CELULA
.ic v(q2)= supply
.ic v(q2b)= 0

* RESULTADOS

.tran 0.01ns '4*period'

.measure tran Escrita_0 trig v(wl) val='supply/2' rise=1 targ v(q2) val='supply/2' fall=1

.measure tran Leitura_0 trig v(wl) val='supply/2' rise=2 targ v(blb) val='supply*0.5' rise=2

.measure tran Escrita_1 trig v(wl) val='supply/2'  rise=3 targ v(q2) val='supply/2' rise=1

.measure tran Leitura_1 trig v(wl) val='supply/2'  rise=4 targ v(bl) val='supply*0.5' rise=2

.measure tran Energia_vdd INTEG i(Vvdd) from=0 to='4*period'

.end
